-- ALU:
-- Implement the ALU using the 16-bit adder, 16-bit multiplier, 16-bit multiplexer, and gates.