-- 16-bit Multiplexer:
-- Implement a 16-bit multiplexer using gates.