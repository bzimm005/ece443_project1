-- Full Adder:
-- Implement a full adder using half adders and gates. 