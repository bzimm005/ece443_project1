-- sixteen bit adder TB