-- 16-bit Subtractor:
-- Implement a 16-bit subtractor using the 16-bit adder and gates.