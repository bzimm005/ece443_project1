-- Implement a 16-bit multiplexer using gates (structural model)