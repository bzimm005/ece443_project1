-- 16-bit Adder
-- Implement a 16-bit adder using full adders and gates.	